/******************************************************************************
AXI Lite 16550 Compatible Uart

#Included modules
The modules are listed in order they appear
+ uart1655_axil_tickgen
******************************************************************************/

/******************************************************************************
uart1655_axil_tickgen

#Description
The tickgen module generates the timing reference for the transmitter.
By looping back the external port, the internal tickgen can also be used
as receiver timing reference. The tick output is generated by
dividing the clk signal by the value of presc. Important to note is
that the tick clock has a duty cycle 1/[presc-1]. The signal is only
high for one cycle of the clk signal.

#Port List
+ presc [15:0] unsigned int -- prescaler for tick signal
+ tick         bool         -- divided clock signal
+ clk          bool         -- system clock
+ reset_n      bool         -- system reset
******************************************************************************/

module uart1655_axil_tickgen (
    input   wire    [15:0]     presc,
    output  wire               tick,
    input   wire               clk,
    input   wire               reset_n
);

reg     [15:0]     presc_r;
wire               passthrough = (presc == 16'b1);
wire               stop        = (presc == 16'b0);

always @ (posedge clk, negedge reset_n)
begin
    if( !reset_n || passthrough || stop ) begin
        presc_r <= 0;
    end
    else begin
        presc_r <= (presc_r == 0) ? presc-1 : presc_r-1;
    end
end

assign tick = passthrough ? clk : (presc_r == 0);

endmodule

/******************************************************************************
uart1655_axil_fifo
#Description
#Port List
******************************************************************************/

module uart1655_axil_fifo(
    input   wire            regmode,
    input   wire    [7:0]   idata,
    input   wire            write,
    output  wire    [7:0]   odata,
    input   wire            read,
    output  wire    [4:0]   elems,
    output  wire            empty,
    output  wire            full,
    output  reg             oeflag,
    input   wire            clear_flag,
    input   wire            clk,
    input   wire            reset_n
);
//==Local parameters
localparam WIDTH = 8;
localparam DEPTH = 16;

//==Signals and Registers
reg     [WIDTH-1:0]     mem [0:DEPTH-1];
reg     [4:0]           elems_r;
reg     [3:0]           wptr;
reg     [3:0]           rptr;
wire                    valid_write;
wire                    valid_read;
reg                     reg_full;

//==Sequention logic
always @ (posedge clk, negedge reset_n)
begin
    if( !reset_n || regmode ) begin
        elems_r <= 5'b0;
    end
    else begin
        case( {valid_read, valid_write} )
            2'b01:
                elems_r <= elems_r + 1'b1;
            2'b10:
                elems_r <= elems_r - 1'b1;
            default:
                elems_r <= elems_r;
        endcase
    end
end

always @ (posedge clk, negedge reset_n)
begin
    if( !reset_n || regmode ) begin
        wptr <= 0;
    end
    else begin
        if( valid_write ) begin
            wptr <= wptr + 1'b1;
        end
    end
end

always @ (posedge clk)
begin
    if( valid_write ) begin
        mem[wptr] <= idata;
    end
end

always @ (posedge clk, negedge reset_n)
begin
    if( !reset_n || regmode ) begin
        rptr <= 0;
    end
    else begin
        if( valid_read ) begin
            rptr <= rptr + 1'b1;
        end
    end
end

always @ (posedge clk, negedge reset_n)
begin
    if( !reset_n ) begin
        oeflag <= 0;
    end
    else begin
        if( oeflag ) begin
            oeflag <= clear_flag ? (write & full) : 1'b1;
        end
        else begin
            oeflag <= write & full;
        end
    end
end

always @ (posedge clk, negedge reset_n)
begin
    if( !reset_n ) begin
        reg_full <= 1'b0;
    end
    else begin
        if( reg_full ) begin
            reg_full <= read ? write : 1'b1;
        end
        else begin
            reg_full <= write;
        end
    end
end

//==Static assignements
assign elems = elems_r;
assign empty = (elems_r == 0);
assign full = (elems_r == 16);
assign valid_read = (read & !empty);
assign valid_write = (write & !full);
assign odata = mem[rptr];

endmodule
